-- megafunction wizard: %FIR II v16.0%
-- GENERATION: XML
-- FIR_90TAPS.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FIR_90TAPS is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(14 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(40 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity FIR_90TAPS;

architecture rtl of FIR_90TAPS is
	component FIR_90TAPS_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(40 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component FIR_90TAPS_0002;

begin

	fir_90taps_inst : component FIR_90TAPS_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of FIR_90TAPS
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="16.0" >
-- Retrieval info: 	<generic name="filterType" value="single" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="1" />
-- Retrieval info: 	<generic name="symmetryMode" value="sym" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="1" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="clockRate" value="100" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="inputRate" value="100" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="read_write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
-- Retrieval info: 	<generic name="speedGrade" value="fast" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="reconfigurable" value="false" />
-- Retrieval info: 	<generic name="num_modes" value="2" />
-- Retrieval info: 	<generic name="reconfigurable_list" value="0" />
-- Retrieval info: 	<generic name="MODE_STRING" value="None Set" />
-- Retrieval info: 	<generic name="channelModes" value="0,1,2,3" />
-- Retrieval info: 	<generic name="inputType" value="int" />
-- Retrieval info: 	<generic name="inputBitWidth" value="15" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="-0.0011117461774144577,-0.0029434772937896154,-0.0036799190313550763,-0.003011534572258722,-0.001163757694486502,0.0011775299748945898,0.0031197334191662308,0.003902944427194778,0.0031962912944831917,0.0012360407811005576,-0.0012515884638817118,-0.003318442554144962,-0.0041547472934654085,-0.0034051992222271826,-0.0013178977864714701,0.0013355876896455699,0.003544186945583385,0.004441281589566471,0.0036433250419633588,0.001411365714589999,-0.0014316731349438272,-0.0038028867226332767,-0.0047702654110158395,-0.003917259255644805,-0.0015191035553984132,0.001542655548505347,0.004102326622053209,0.005151886643897107,0.0042357356178923606,0.0016446493037784301,-0.0016722904685478306,-0.004452952829066315,-0.0055998767868446825,-0.0046105794778828245,-0.0017928159077224533,0.0018257116124512807,0.004869116644866891,0.006133198385591793,0.005058208553405442,0.001970322433239528,-0.0020101269268402978,-0.005371087432997514,-0.006778798215654088,-0.005602101946244723,-0.002186841381947122,0.0022359838849122407,0.005988453804606422,0.007576303888083979,0.006277053987960955,0.002456821799471459,-0.002519019819711258,-0.00676617507793193,-0.008586477739828511,-0.007136924397270675,-0.0028028530388336677,0.002884095155901294,0.007776051955235203,0.009907474315186742,0.008269769539694593,0.0032623371435605,-0.0033729248433421897,-0.009140271596504537,-0.011708833281584334,-0.00983010341510867,-0.003902011093278246,0.004061276852187533,0.011085010234058707,0.01431079623304752,0.012116173976761834,0.00485372111602904,-0.005102629891209976,-0.014080958945966464,-0.018399595156775382,-0.01578774184850785,-0.006419437605070633,0.006862157439903067,0.019296128925954042,0.025759433219485536,0.022651977434815618,0.009476312655104272,-0.01047381925037842,-0.030646793000044626,-0.04293238869914256,-0.04007657546159684,-0.01809114234156273,0.022111396195243323,0.07442792585725129,0.12879716609742767,0.17366516033358634,0.19900256575718986,0.19900256575718986,0.17366516033358634,0.12879716609742767,0.07442792585725129,0.022111396195243323,-0.01809114234156273,-0.04007657546159684,-0.04293238869914256,-0.030646793000044626,-0.01047381925037842,0.009476312655104272,0.022651977434815618,0.025759433219485536,0.019296128925954042,0.006862157439903067,-0.006419437605070633,-0.01578774184850785,-0.018399595156775382,-0.014080958945966464,-0.005102629891209976,0.00485372111602904,0.012116173976761834,0.01431079623304752,0.011085010234058707,0.004061276852187533,-0.003902011093278246,-0.00983010341510867,-0.011708833281584334,-0.009140271596504537,-0.0033729248433421897,0.0032623371435605,0.008269769539694593,0.009907474315186742,0.007776051955235203,0.002884095155901294,-0.0028028530388336677,-0.007136924397270675,-0.008586477739828511,-0.00676617507793193,-0.002519019819711258,0.002456821799471459,0.006277053987960955,0.007576303888083979,0.005988453804606422,0.0022359838849122407,-0.002186841381947122,-0.005602101946244723,-0.006778798215654088,-0.005371087432997514,-0.0020101269268402978,0.001970322433239528,0.005058208553405442,0.006133198385591793,0.004869116644866891,0.0018257116124512807,-0.0017928159077224533,-0.0046105794778828245,-0.0055998767868446825,-0.004452952829066315,-0.0016722904685478306,0.0016446493037784301,0.0042357356178923606,0.005151886643897107,0.004102326622053209,0.001542655548505347,-0.0015191035553984132,-0.003917259255644805,-0.0047702654110158395,-0.0038028867226332767,-0.0014316731349438272,0.001411365714589999,0.0036433250419633588,0.004441281589566471,0.003544186945583385,0.0013355876896455699,-0.0013178977864714701,-0.0034051992222271826,-0.0041547472934654085,-0.003318442554144962,-0.0012515884638817118,0.0012360407811005576,0.0031962912944831917,0.003902944427194778,0.0031197334191662308,0.0011775299748945898,-0.001163757694486502,-0.003011534572258722,-0.0036799190313550763,-0.0029434772937896154,-0.0011117461774144577" />
-- Retrieval info: 	<generic name="coeffSetRealValueImag" value="0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, -0.0530093, -0.04498, 0.0, 0.0749693, 0.159034, 0.224907, 0.249809, 0.224907, 0.159034, 0.0749693, 0.0, -0.04498, -0.0530093, -0.0321283, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0" />
-- Retrieval info: 	<generic name="coeffScaling" value="auto" />
-- Retrieval info: 	<generic name="coeffType" value="int" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="18" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffComplex" value="false" />
-- Retrieval info: 	<generic name="karatsuba" value="false" />
-- Retrieval info: 	<generic name="outType" value="int" />
-- Retrieval info: 	<generic name="outMSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="trunc" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="0" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
