`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QuXJLuIQ9UUx1N65MC2rLe39xvUfYKlSujjyy3aNHztrpA6mK6YfiOXxQFI9cBwCaXCBgqcYW+B1
UAzGGL2Scw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SkqHO/Qm/mygFtINmM3LX/z7CSTLycUvwRtfru5lwBJGcjg0GdHV4ky7uGxR9eQs14l3yM6a7alu
g5jXxGp9994dzQyURFFGUiSNbjSCsAxIfYML/ThEdVv0B7Y1PkdvyBRCgTr75Vu/BYO0+BjpFsDj
vsx/9/hY1XS3ZYi25CI=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V6eQuN5kCBnirWb7KEYAe77sYMrzlxkaawy7JS9Lg1qGC75EKFX4nth6ewfwxAwFR0VQhr6N87vw
eW4yOHwE0t4d9oPW2Oegy/W3JRGIQQ3AWo3qcHYag2gXzRcJmhLV15B91AKBp4czyDtXcSbZYCE/
JbK2m8fdCAZGNPFi/Ao=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JC+fCbFN4J5J+65rf+U2mv0kAGlqfguyTeFXZYaCFRtv+HUST8VWJHFt+VKA1jqOTQY2BSKfpEZA
aRKhrIaZedpTS2rA9Ovr/0mFCacHl/jeuEJIr04GICikqj+74dR0lsCkoAKkGRxYZgWStJTyRYw9
H6miHw9Y1KAhXMBdNrq5BkxVPG+1cCMsORT5SHhB0eAWKL5PHdEYbOgKWFu2ElsKE9d3Vg5R11Wi
Eraf4Tzqg7ys0DtI/nSEvdAaHwK0OB3W5YFjALNdX7aOWTIyH8AiJdEadERK1NknMpswiafPpANT
V2a1EpxQ4oMedAJSdIW5TmzdNvAwQ5dY6x1mjg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bkk8YDXwb7MZPWUI37XJK/SeR0r5xbQAsT9ya5Q1NIsxqHe7ZM5ve0ZAuBhb6QJ+fIBHB3FnI/SZ
aGT7YDsQhpWPtcgs7EQ2dK/6qzaDsSmc+1H3iL/h5mlvvmgBv6o8Tn/jYJpKmWwPRC3GT+aepkyr
eoERGK9rxvUbdN3qUXbVtyRTrsqgXNjDw3Tcivjt9dSlNNuQisYf8h4Xi8czhv5E3tX5WY0lFIRn
pAPMt4bMH6LCe7p2XrWkD5S09+1eyCCp+2EOwluC4LJRklBR3R2C8Zk+OFZ5YVgWgoa0Hq7+1yeW
XHikW/W4VFz8A/xVR7nb6Bu8sByJv/YGXealmQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ka1fgPqQFifFE9IP3cUwtR44Wg4Eo470Qn/Lil0X4nqk2aSIMupgwScLReHRc/S2+wq9uNQlBhW8
cRfvvrXJtp7E9hmZFKNZUSPqQIOWWeDzXRLnJ0YQaW0V8zZA9JvsVkdKBBtIZ/ZWlsKr4i/Lpqxf
Ekj/m6a2pAaevsEeCg7FwX/x6MX2UlK5/NLka1zKjWuUz6U+T2Z3YKz7nf60+YFJLQD3hGno0IDH
wTZExwOd2jezNdQNM0o4nxcpAywqXOQWD04rDfPJJd0AvWTHxbi5782EuttqZHENLv2PRsnP6h45
NW5UxVO4J6zt/5g0JIumpHHyQNTDXgsuWHE2RQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12640)
`protect data_block
e9kUx6L2fEDMplH/J0Nurgy5svvp0m8ZykizEoz79EyyWMO9E1XiZT5Dkgse3D3GqCu2V7zEtqE1
mbt5qg+HUh/zn0DPidgPhxo5PgT6rqTR4uo+i1AtPg7xjZ5/wPqXsZMiw2B2nPYKXFYo4O2fGaWc
GX0kuV9IcyqafsCVqoNLNhhmz5sqjkuHuM2UetSXKGXP61Dz/6GVtg8q3vFIwh1vmOjsP8GsxxHe
ZZVbacrcF069HIBhev/E3frgFH18I2BRCnIR8v7pJMetPuORzekGelCXLO3ot7gPnZ2e34DOxOfZ
4wZOOqV9+EGPlMNCgIwgWn/MZBqtUh5atZ1VuNjjRQfwwFkoxaXxOLwDkj1uf0ztBxLS0uMovv23
s1fIzi1ORAS1juq2OdEBs2onY0NiLeI3pw2LJ81n1WltJbMRczJ5xx77jg6LHjuyRFq50EYFCcx0
AFor5xbvzUPPkZZLf3iSgdzxsXVuQnsTeHwrAsDuQAkDHlP0wsiMV59ghf+8j+3v67j8UpzLQoOg
6nYQUFWUjUiuMwCODfUN7SZ54w2igXmbnreIWs5G/8cjDSEs38tMumlLJJ+S261jz70hX+D1Ih6n
XvYc9exey+ORE+etpKZ5LT6n1HhRe6APYp7fHpAy1TyU4SP/2dk70sKrPgIAZSEz2qtI0zL8Q5Hs
VOIMc+SkZ/CeUq9eC6lj3WkfgvGy3QztaxyK90bSZrtxCd3zzUom9omYItivihy3EQciiQi8MSUB
mWEZXgmgk6jXaCCoftkXd3jM7YhQYqAThQb8J4O9+gbyld+zKUcOKEBKK6FvWtsOgZFTZ2jZZOQz
TTdZiam4MOpXPAwtgJVeXZaJbYJukl5y9YclibM/BLQH4/mcISEDRqK2cTvVy+6P8znEJEs40xxi
xK2zd38lDsWbL5lcajeS8VNSMrwl2cV20prJZ/TZljsHnblNq/+5pgyf/2pwHloPqwwmzdqVdzDP
3/x/Aso2zF0ODrlIIreK9/YoKzsjo6c/Y7q+vCR+PgF2Cv/HCua1KkyY02LjFUR8aVMQjc4TJtEg
nAgpEOjmxle/O4AOqHUjPXYqF6mmlMqApuAmQLxYTMt3bW39Qsu5wlYvIjbE3eJ+0DEgk6PC4vSZ
umlWu1KAp0H2ljriaTCF4RoB/ADo/uTq7f7Jedz6rscVIdzSjQhi95tvSpipI8xHyOXNHbxQGqyh
JQMJbsrpiJjoJfwR3AHvtCUfMNYk0i6+cwSm1JjNdNFjBi4LJCv7OfNy8YBf/C4Mr8Ywt6Ij34c+
EKYb/DYNIR8EDhDtfrgvBx3Yh9U3T9gaccfjIo5IeyM+TcxshGCNjKbHcbFlCMyfv2aeByXjjYu1
P9q1uoophPXQRW5Lv2b9KtAz+zre9DTcmofRPp7l1mwwPb4e8S3C3/TgBpyRBoGq2gfMWxhKKqAB
BOiRP9YA1PvAIG9HvbumLxFvzxFTuNa4kpAuZT9kyQ0sQleUOZZhHi4O4n/IVo6FUAz8nG00PSPG
1KBLskjlDeU3PSjCtmPUgf+fdliWI1pt97ImbdtEol8Ex4Pzzf73stf1TfZyTUyOoorr0HyjV8yy
iNF6h9TKlvKmGimp/pV2PLsbcw7zuS0iId2SMrp7WtZ1rOtY9DJKqOSKhp5kKCxyBDuTFjhdBEHB
qhaiXyqQhFeM0b8/KAZui3UHHecZ+r+/1tW1U4QRzpayBc6Z0bESC8MnKtYjY6H6LBvdT1BhyX9r
NgUIiM6LquSmUtM3mWr9EfNRgJPTSujFWFy/tnhUk4pY9AdGREwIBgKdLMUtCM0ku+b++1qGmyLn
LSgqmi/P38degMxQkS220+qrqKN/P6Haiz4PolfDztc5xV2TBnvu0wZKIoIh8San/fAl1kziOhnM
fi5vRG3KreNCkSixyWgUAFhw8SohetGCD1T+vZ78u4126t2xtLW7kXnfILAMPEma6P6L+AaJ1BkU
M5S/eBpoAYVfi+nnr+IM9yh5mdNn7XMXFUmCWMvv3yUW4kmayUyz0EEs5H+CTY/U3z/HwZN8kljm
ms3zi87MLvDi2Rkk3L/sopJqbqHOQZ8/RreeUp+qZf6vZbgQEzAraZeoXOts3TrRoOyUSSgI52AC
PZFTDnTiLmm5SVaAqhpikZsCHDE+GrcA8QkfTdToTZ4OpV2EJfZNtTXXxdpIea7LDZVISl7nMkza
Y65iYl0OTAjIb8Dw13jVHUSlO1/1C+3qMOCdFjEqXP9TM/gP4HtH3AIDlV0HdgbIz51bvFpmycDh
FJQWwH8JCelI/0zKkf0O0CC3Xw9MrqjdoNDaCipY2hSne3M8TqI/7qPghJJe7Hy9cv5vCSFyYJ2v
V6rhJB901LvU+CmEJn6fjJFezDzfmaTdT03gwY7dXOfb91Ex2gMWh7vIuiMZPnoP8FhRDs/peq+J
MptJBlEWZ5LyofeyXgyz4sEwsli3RIsOc+efsDejVWSH/Udt3M8N8csX9IE39BHe5MDU7Xbi9+S3
XP9LLm+gAQWjJXyb1BNVCBLAIxPvx3ACztv2ZgPCzV2PAvqkmoHUDdct/qScCMDq605LGRjpDu6o
k28YJKGWNYV57TMgobQ2lzu0RY+unSeBiSIoupiDiSQaiXrJZD+oyh15uVJAdCiSsLdp7JaTCiZj
7vr5h3mT7r5BOECdSynlGnzF1XBArGMEQsB5sBg6BvA3yt9gefAGtF4+smUnzfSHstsMiYOJYbMv
lxQHUPjmWxdMIypEtIPnIqNUlKMNLv7YKN+l03CMeBJuCHnTnzhNF2rSVfuapysCQ3x+dw5nmra5
0fzFIG3dXClJ0AcPRhUgOdBSKHuKqTeOO09iZAT+FwSVCVlQqFa2JUO6cXDjzxDA/yR25id21gb0
ICIuNeU8o/rAVNHTj1HMjfco54q/60FIVQRNXP/3vUFoJUBFlCdToJZYIac6+6rFVtPCl6WEhFLm
GvqhaxrAbJy2X4loOPbwITtZDF88M11s/is+RntxFFprzk5Sq6FGB+hG0Ai6ZQJhEjI5IloJwBjh
b0Cq164Xq+bI1hRNIaDbLeYmkK1gNUYyIJzXg/WLGQe7hhNJuOod6shVSXMLu9G/JUTpe/wsNCJC
y6w60Kok46lUC02o/bbsiv+VLj3drF5SQuFBSrqzP5ukNKjXXoTHJh7i5fUpDlF/gxKrZFlQzwlh
kV3PIx96m0eENE6SnEO0lg9XsngD86KxAVXzEy7NXJ0C+91NeTI+ZCp5Wu3PLHIHhgg2PmT6w4Wp
WfLbwtVW8TBRMxZg5WvzTYgZ6tov712dS97seIP8MEZ3dHUGCdfSPFSLMYBiirvgH8kggz32Bn1R
JtzXHCmZOy3owKno0kGEJrAQsegdSm2XTS7jQ+o8FlR9181B+HeoQKwBbmFEkuhQSOA2tRRplxne
sa/SdHE2lkdJLzZ1I87s0zkIZwTZXn4OaPox7pBRGyCUYXqC1+JgUBwdcM1QlWN3U5UGGkJlOv1z
0XBzPswQ5Iu0zQBk/Leea1I5S6rgM6/kyuHSzDqKywwPCSsa04sEF2zLVpA3/yy6EejP7pbA9u2l
LsKa8RDTfUsnUEjvUuh1vc4TYXmmTlCNKi6oK9YxXFj9PYKvSkxMh8zAF0aC6/3COyur2CtsZ8mZ
VvVGMfVXEuzF5dd0ZKy6MZFF5LGH49gsjvKECqpPjmbipng6DC7hqoBwaHX+v0VBYiXXoG63wuJM
nc85BsfrbeFpGuVNFprgHfEle6ROHXVgg27U3aW3fZyNdVMnUSugRCbXXqgSlPYQCAeeer125v95
VwIrL70bySJigQ6gplgDiSh1ONMOvRkIU5PEHuoLOX5vo6hWoYCoIWMQ7lD5rQAP9wghYa9xTkKF
NxRBrXWOmG6/B71xEHwHas+If14QMmwI+Y+ifxpxTLa/vAoASWUG54ek/kRqR06egKHHA1WSWLBS
TLQXHqfKQ4CMARxArFlT22HXMxxV0wCqGZ855gyOYQOQBhaNYpSbH2vS18IeeRNp2jTSQTz8d9Dw
SEAxT4iDrmUlauj9ETbTCY/R+sAZhB0uU1yMkonD0FprEtzbFD/GrZPOhZsAqMqqxekL9lycuDLS
xFeedt9kTKf4T9NkMt4R5xd03aDszFcm9iCKmIt6VoMrG1enDhbIo3wlpKBUtMD+QMgq37NgP7Bw
SRmApjB/IwxXv3GtgjJIzDSxiOErKtw5JUdRffoIXz8yxjPM7rLMvVGdZ+fCVJ5N2+9Xrrt8Upfk
hGq79OVmEaKfcaxw8RPLSKPWNlFBvnpy5YiI10dJ+uCcul0b6H5+0LvCD7CF94/0S9d0usPctrwA
bBA+NNbLPcDLkgG2/y+e5C7SJ5ryeaLjcC2mSv0s+pIytG7zyp+w2HHWWLKvH2hSIL61FZRCa290
aVNAdJR2QJpCAbv0aP6MHsqb19+dkMv03FaGGfvElkHFh8bOz65s9dzEM+86SAsRh5PTlJ/NDVO8
JsRWWVd0nhDExmclGgUl81aAQNaLsJZ6LHTWlaSj71+ktjddBtOCM/ljaBaSQ43FIsodkAZfPTUB
QQk6rQxPoRJWaDKZfOqJKR+gm5PyjLlenOM8hGNYRS6CQeXtYyFriu+GjPwLFdXyJLI0btf3TCnm
P/GqNqjTjDgGggXgNxTbJoI78oIcAvI4hf5D0KCT5abgefO/cy1RrUF1x0UTt4VaCKQjyCVBpOdb
eq/hZrQbobLeLDk4bVk6YR8VQojaBrZmdgXt2P/YZWhbTbdgfA3q/eQWg4IvAp0KnxLAOzFuOOHO
qME4W/G7N+BMFV6SuRjifg+0kDdIT9Qw6+k+jqvBcsAOP+j7Tk7IBvzaPeE/UQ4dQsa4uEpbLC+Q
bTPllDz1Dt6Fs+pmGd+vAWaVTr4fKRRYLq7hwYh5892gFNK8djZF07G3K1NW7ko1yfBw5tmDkado
6le836TPpMV7pG9/JchMvVunIi42X3JAWdjHYJYUJ6ep0rC8stzK7oHUZGMCTRYsE/7cL9A4HyV/
vYcP4zhTyP0DguzHauhjiJgeuMrWcxAfD0nX6MgbdMBerjRiSoz6XO3+PzPrZ+SvIhrqCQHVW0Xf
izeO1BTx+SnIkG+MsYiMjDSdZj2UnmeB63ilDBILqwqbg8+Ks5JucsX/SEkR7yVjK6x7nLBcKe4r
B5ktSmHFfy5XIafrrpLmTR/zEm79TO/wa5OBDxiWOyoXj6kt0aPfZJDg8I5ERpTOkmX3vpzTYrOY
Y7CfkVUVgRZuopB1ToI+si7jzsu5HP9CqROogJVlN9RPGvPJ3g28TROAabLb+DebMfMZwEqwXyP5
v3/ujSJfv8//iB8XSK/Ojy/diSNLki/zKjWWUbWMXq0gQHqr8gEmaydF1Eh4ePyqhgij1cd6xPn5
dlv1mANqmHtYELoNLTR16sYkyn+TkdlmqPaXmX7MuPNS9B4t7t/9rDyRCFrzCFq0obqL2qcvtWke
LlVFH3Os3ocpdrZvqhYI6Rw6UazQ4p863VgweYJOeB+mGqiLIDJykFZWMBdMhVutV9gQLRICn8o0
qujim1lyoxulfjm5YtFN1CrPEjplqkcl+YsJVSrSeZBwWF8SSdS9a//WPZxlRPYxbGcdQw9439XZ
Zk7nZAzVAYvM6toykx30Z7G9mPdsQeFPqE+nY2LHqxYcY/5IXgQf6Ndhd2DEf+BCVzgOXQsuKtDu
eNuDgv7uJsCADoP7J3mth67rOA0qEnah0zWyb3ly0hSoRHaMZD0hzzx9rSzP4E1O3tSDIKMDKZHr
bsFOP0NxXO+dFjB94PSuLpgfSlRpbWHMTekh/mIP8nk26X+6v1LmGvq+3lpwjjhA1AK72VSTPDnz
XI5dR+A8y8/ZN+gRhDTP7ia3kVuGMfol9/TYZD2uAARpR3LgP35ugiLcAC4j+yNHdeYKVpXbA2uA
R03Lfkw5BjPo93ZQPckjfsB6CNuqC5jGvZYVDQ7oOyz+owWlRpMr+j7B7b9AN3xB2GWFbu7WBKLd
eJfF7HMRrNbRdnBiWxFC1w0ryHDTQNdUUXRnSRU127HiVuavhWNIGDvL2rhMHF8RxDvszYA6Gsie
oW+YtcmntZHyfFld9eUsEXqAAHwtsMDYGm0nUPVaMBrTgbqHQOSSePGlsjD7VRrgKnVHF2UYgqee
L5UnfB6vDE2dGAV63Y++nvEAnt6Se8Z/6yOwjk3m+MZzbowVKFUmDv6Q74Gd76ENr+OnjzomV/tB
/FevprZSzNPhi1OMPbmwZXDdNaeb3gClr0o+NCKp/rUGPtozHY1ijJbo4jZ/SHPZyFTtU9oLkrI+
zaFSl7PEMQkEqLx7yE71e0jlGeq2kI2tkccMfWFMrXDV15cifkz+f/uTw3bQP4pmxrbebzZpDgCa
CXemqqGjwokv9KtnfHRBfGmZ+wnXAERk7SfyNZsbcuJiOjuI/Kf6zJYXWIQPRvk7FGJmFICUY2kG
pDBq3PRh9T865RTINE8ngyfIWz4U0qWd5hUbDyeOrtVwHQhINQnM1ZtUuMPNsJCHE7IR/AjAhKEh
aIokL2H7IniVYPzCPDOrQ1ZYs7j0EBgZ9fCdPTin3K4dr7eorl3Yz4RqcaC9+tYnBg9bYhc0KFU2
GsOmW6NmF6vWiH+o5n8zMWoBhHs6A/TctWWlMiGqM7wmM84DmN3OGRwMIBspMCuENQrAT7Xw8QhZ
AIVBftsyLtu3Obc6aeZzXwrylTYAPWAUjxq2I/MFwE/yz7ZZd+td92pEBuUBirURcGyNBMBwJScl
Ja5j+oW6YAG2UYHpiDPM30MVH/mHj7nYNUvwQTas9ER9U2dz54y8zmuspdphFn2LwbhB8CbhcTVV
n5NFsz5fEJt2UIXvDGAMFBNAyhoyjrqQx97TOm3w3Mv0CK/bQMjHl2cqn1A/3/j+V3K0SW4D0NJl
LOD8JDq+/Ip9u3HtfpzzQ+JWSSUo03f7YLmnee9IsHwNy0EcoYuGRPLuUcc0iJVddUzxdmKwCpnb
8RLpykSl8Vpbyub4YuOdnz8N1nWfubjJ70ibpA+H4Rn1JjenOn1z475zNSsk+uDvNO9QGHbu4cJq
CxJ0nWcec7VhpXgcYAMCM9DZipkpHnGYjlK8dnCpwGbbryaGB3UJgO/d0laDNuhycn+vqxeSmPZD
EP2a7dlLG5OpBmchiTPhn8JftyH2dDZeM9eWsUbglXTRrtj3xaxI/AAP5xncQjUo4ygPlnfw5sze
C9j5U9LZl4n2CIiiCFWQLNVAD8WKFBSBzdacNH/bVTCsf9r+ECbm6z6Sfqw1X7KJKXrLxLcskX4t
xtVKidRjTWslPq3azlsGk2sx/dctSjN8Ar4sqLgOjDnOAtefWTHBiSwIA3K8S+6qSs0E1a+Pbur6
UTytfoWIjCmGqX/d3Ti70Ic1VRYvF4wYuzWuUVpvkN+ipvBVN0XuNNIz+ftU/w3Yl/VvLDORkTx/
i1D8C8wa1PtcsUQdQ5ua+OIhkNqFzd1ishNSfVlgks69WeqAE7jXOlPrOUOaOJuzvFAocLgko/hd
Hr1P16CVIQ40AvUkicO7mdeAHyRuAWkrEoxzyVFI07I4vyZqUjDxauvaNez7aAqySIWsh7Fw9XKF
UsRHlRBrmPEJK48QhsNGqXJ6x0Ht/v0BnzUHHBBNR1/KddWPfcLCghg/0uPIcJeP82kV26JiSuzH
ke2EXlT/QqBc9wZ8e4IdWMZn66g9nRymVbSBORI7hglYmDpbGL7pONM4tYkaPBP73FP9eYXD9AYM
0ZnfGqbW6+GYx5IIgVi0vqKtYyczpN/2KfUKxHs/gP6rHn4B9PBwNjk5uJ7zpCl7CH1fjHer3qlK
DqDlTXWyhFGFP8cqWGeLxcfZeeTcMFq4TNbDzJJC/IAvo9K7bSuXrH/coKqvsCpS3VK+PiK1fL52
hBUVogN79AjUP7yd6JiSaD7MA9d3HbL5N5lZJkPjflNtTwdk6pN+jXGrsn9X0jbmTmsCbYrKmbeP
82cgPMRKW4XZbQHS9UteeAZy/0SlzeU25BUYW7sSrU7LgGvyWv6qmha89DYnSEPKlymSp7wCUc9u
g4W33p0bW76EtG633yY7mT6M22JMQdJAhImHfsdTeighjjXZDaEkHCkoze31iGiozHhQP1eyEFSe
EkkXaRgfHxhl5R206hgYtcVX/aPkqhfOUZWDVUVa32NfBIa/uGEmQ1AWgQorbe/SQOM3ufQHFsjo
mb+w/TMS+mwa8f9T+MalikNA8XVBs7moW6GeNI2qfL5gOX14JW4XSjG5+ejxKQOXySjfgBeDF0ig
zCPkTUpjI8Ve+6kub2hL26REbKm8QtgVf4/Tkb4+WyKz1z5kbql+4UV7KZEN8izowDgdWmJovkto
xlT+1tWQENFkCwklGSRqgEq9cFif4p4Zzt7nZa+d45UGKSRkhoVCdaOlfIitRKrSDh95r0OuR7fC
pTIOwgXCncUbopYXCj9L2rpTYmQlrKA85dZKZrQ0oZaOR7VGlSidgV4Jtdyo5j8hWXRc7oJHUGfI
e1SG6skxx6oqhCB/HjU4Rm0dwitw42FbE5YpN14+EvoGvmpj2BSZR6yruTLlRI/gpC6hv6BvSp5T
ZGajrIgMrbsDZpv/G0Ww/Zlz4bw93Dwhowb3ElpM0mqfEORY/0HWsLFspHQpk6pcKVcx6IrXn1Zp
06h0VONV7dGVMppmlC0y6Qum9ppOPUFMBaYt8CmkyD+uMmjrOZ7o4AK5ASaao2rtOC/GVeqemMfe
abmS4+35h/PkRvmUYrE+WH3KDxGdCUO/cTh+47AtwwIOZ0BxajtMeiiR7fXS8leeLXkAWo0elEdu
lD1mYYeSV+MGcLtyhMz395DQqdAQj0OxglKySigNqLJ+b9HrgDBLLHo2NbIQ81bdswgHiSgGiYK/
O9I62Kvq42yO48gD0HkLiVcGCfQfWnMncMf/kGI2k+KqRwcW0cZkzyNfzihBuAx2pDfXR2gfs5JM
I1Aa5kXlfcxe3mURDPITHub2jFcSCKeKhaJPo5J6UxYR8hiPz3U5QJourB06+qfReLi+Rqt5EvxF
gHvHBMhS0/4fc1oMyzU99mcWUeuDsf4qJS2ON3pmoNRTigVxYSa7F8WzrsZt0uBwGhDNuu41I0Wd
NmYcQz0wsfnUIdbQ6u7Wo9TBvON3Sqc01DyFSyLRA7RorysoM0GwRQ1uekFFDr0qhlcZPKp5GjHk
d0PIF0y7sNJJVOHets8v/ivLntdZbLO0SvJltbQW1BZkAlAzdy8EfPGYN888X2kcE+zwvmVkBXNF
QH9YL7NwHG7Diiqpg7lKwE4pSNbdZT4t6NTF4PfGdLw45K6UT4mdccPr7qSgbRMaawDdvdOxVpk8
JvSlR0bqMISbkNjaEujmgdjccfm+uVgZlU9mO8DRtlpWRVkTOG+mt2+sye21blO5fGk2r70HeCMW
AWjD+9JingPZFRS9PW+caTduN4w8wjDj6+t3yYGkl7Jnyt/dEseX2HfaaGlHN9sybKMc06+oGjM/
BYDle3lXwf3RadfhrKGGGARUCEfutueff9DL9A91rhkYrKkbyVUqQRgs7tG0W4nlNs0dXqO2ZDHj
GyT2VZaX+q46rZ/0vhxjs/J3WkCQH7QWO/wtKUBCQpQTlvUH5VFtl3gcOIJn6i70QYaLjSo0DlG6
BQByIhqoRObbv7f7jgHBdMSu4wh8pItpMK917g0D/2VBaQoEuJyssbF7mpR4yr0CR4CkfUVa6WkR
JHYv/0MVQnGXsgGF48jlQ/5bY9+ALEV9qJvE6il5DkgS25BcsAg58MgA8IWw3JViGZPCBNZnDvi4
8+ThdKdGVjb/1dFo2U1gQiww+nkwQOOET8jat4hIK3fn1Wycw4brpz9a8My1tZNhpoG23MR+cnYC
tzrz7lihiYFNgHlm4dxAhMOiQqSjN+k+tv03qFX7v0BT2MW+DaQtwrooxj9l4u38wAl9Y83ZJn5K
WdvT2RDVHkH8yOHcxLhwtFDyTnHBgvtDZ7L7qr6zoELdLPbYFbTeFImSP2yEt7LH0u4qxlf8BKO+
1P0A/AvuPhdTI1ywgqnjNkAFo0dxdDHoDLnTX77dj5TD+/xrnHXW8Z9vOb+l9Ou7miD830LwsxGo
EPtBlMb+bOGsdogbpoecPUxuy6/7UuxP5IsQJnmuBTDwjYV+UpoWewPINDRkwwceLFUx6OxylNJW
iKe3nVpuGng+28DbDI1OGBSMmVCXdf79bHZ437sX77jIiFajNmvWwDYN7Am5DusxYgXNzsZ/lAqu
ZU842gNtvIJZv/mjcYqZMU6XnTNIsh7NamclhgN7QQbPnKd0th0p8L++S+3s54vtBZ+VjkkKcrZL
0u+SFCSfWSgJlJHlZTnYVOFlOkM8gIq+rJVJku98/bfxszC8NyCjewFDetxUDdo2CiNLubxLir82
PIa05nHSBBgdhWL9GuHabAGmWEg3LrmsOyw6cxVoyUhptT/Bx9nhKhWO/JO2eHVEnKuNXcrSxtrf
qDzuTMPX00VY+xWV0NlsTvfgYRfaXedwCEvVWfPVdfmcy4Fw/ueE8c1x/jNlnR6RMfeNgp/94rDU
3DdU1VcHwKWXsqM/lcr/Nn4lvBQm6/VWGgnVpfMdNbBPpHkC03XprvqbSfBgzq4VxyiWvnwVT6bu
fZm7FuFbw3xnVCqA6gQq5MrA/i/zykQNEji3I0OhZwZJGobv4fHZBpvt5KJknFc4NzSNX5eoiPuA
ZUicffQwAklAD7IWuTmn19uLhfYBs6yN421WVHoZJjL9V9OuLK8YwYBMFq22MsRUQT5L2/g9AvNl
ZznEpv00OtKJQ6uL/fTD2wjFdPY6BZ0PX33ksB4utvW/uCWg/kGSKbweT/0ehrOshRvaOslx+vZC
oZLFvffsW7/ELNLwbxVo8f6EIVB2MhY9DJE7UIQVilZ7AD1NLPqCDEp2/C6nlaH3xpMiGWafPWgt
IhmY2ra1vktzHs+eZBtMQonW958ItLFa7KUhnDH0F11S5iRqJ4ewVtQVRn5Oz55tLMDLFznTNv/y
Zz7VzAwgDBRLunMIgBgaU0KodGTn+Y2SJ2PPueqtNGx+Ho03f0znrE6WgtkgnNMdGaqioIvyUn3Z
he9wnj86HZN9218mjrNfvtsEfimKoyZH4Q7qD6rvtc5mK1kTtbMutQlzu0YBXQJ6LZt4caLJacr1
8Jxi8S2JNg1y8hS7gxJiqkWCUB6m6zdlZAJGEeQ2Bnq3nFZ3cdbJK6Go0wnYP5AvyVkRCjTpkEyp
C4Sjg6EDI920MlFIyKYTathnQv9XOoYOqhQpMVD+6MMavLxXJFUhH8jvrkv3Uzm3BzmS+1u2srgF
I5GQUapnJnKdQ3jGtW8x/tlO1D11WLn3Qp4YJ5pDoLsckhppYhx7MI3DFtQPw/HPI/siMjhVCq28
5/nLBnUBP+4dt3VhI7GH2Ya9tGamrDq0FIGJvxPzWzpjJVxUV6LIdTQ3inHBfj1cOUi17mcuPv1h
ui+bNYC2T01N3FHsi/0evtD6nyoeLNhRU1aYU6aQJsnAFxsH/Mg85smTe2iKidG4trynIanrh2RF
Fbc7ybs44go6MCG3T8iZgWTWp+wHtJ/RPg43fCYF+wbpgKQmc8oqUcSZGoDBxsByN1ordx2W+O1u
mdlINvTsPL4hBgzUtkPSHy91cBsGNTEawhJGUVKD3fOfNEOn9aO3MExcrgOyd1mwfLPzaIbxgVEl
FD7lbJiqyfDlFOPyywl+h16jF10BxOff804HEAamsm9Dq15kUI3gInj61L0bVHSsln6Wi1i88DVJ
+1uRSrCcpryXh6Ifgm3+6RtBoGIZbsZYccQC1wBIAPJLnxxPldf21Z2S6kugFwdSEDrbZAS8GScW
OoJ75eoX/FHNYJaprJlJy8lWI2XB6yksWwN235aTaPiErovt4hrgMLZMCoNE9OF2VuNgSrUKUaXi
SQ43l420ai5oYJ9a6DsecvSSTmHDttztZ/LBL90nzUNMTsjgbWXKgurhyQoMSSY+7aGmJJRTeHY+
RabgZ+n71PMRuIAkmkn0PQlsUX8Ta1e7OO21PgXec+bz34rJooTZQlmkhzdhnLRytM6e9tleU1W8
5XOa90bkP9wpv1sB+43yWGkvVYm6zUVEesuYMEbJX9M4ildZDMMudDW5Er+gblOxkjHA46+gh5zE
DRzrzp5aZrR71FaauMCqxK1QbUDCDOSFFqRVUyFuv4W4gbNPF4fHUTB12ztWvOrLB1UpfeYukLG4
urbx/iLE0YqTKjlKgUwQk9ImySlJ/+wrsN5nH7Y6sojEuKt+dd+9JdG0V3fd+cl9oNkrp6cLqbGm
u4yciB58GQG9wDFbqIHL8hqKxv7nY+FbudSRlGmA+MNDsODfWvEyfz3jflaVIfc9aeGbSnLbZzY1
F5HyKzJUI87VFn33TRqGJ6lFjn6z2mHkYWOFxbqpOOJPJ3I9W2LRxlC39kDQ0WQ2MJAzk51lTdWi
t3bVUUX/TzgDNjjMjIR3Qh1xsRPEy5+lXgB/GcEmSKBX7P+GZ0H0d3YnKbU01aR7W1mQLDmCmSL/
8wbGf1XbKSPL1zEt2A4u5HdAYjqkqwQFBomDTRrUPVaGxKWkOAzayCpGt/EWiBw4GX7MyIl70JRZ
62jC/2+0paovVYtHzxZWKDondi29ZNStO1hx6/p4x/M9BKJs010r/UK67FvmKO3ZsjBZ6rulWg1h
MGaDbe7wKb6UavjDcj8sw/7/nxE1rdTrrOZ+ViCs38Q+O4LT7PK8KP28M5KYEZOqFgVWIv1BVmi/
YLCI36hCQL85elGKyXyMlTCGbezfAuWDcya8nAFALNXueyUeHc2WmZ67XJPB6brFqZsoLn47nOmE
wv+mS9Hk35i7FsZXva9FzcS6pgR9PO2IoyZTCQ1U76wwdQxBitJukDJE0FC75YkuNiQxjQlK9jlK
rIBpa6xVkt/4VOAt0hWzbwU4FomnBpaxJnbKHAcrvgIbM1ohSH6psih0ppITLkXuoRaGyxwO6SWu
69OwHCspP6tX1EipEmSc7P6/8mMDotnhv7CHZEvcukLbhpzIQ+rmgVszUTV9k6qv6VYRPOecek0N
KeE7JFFQLSIxoVATVVmLyjTe6ssyNLosigRcxTShy8gO3AWFQv0FYGbf52vSqt11i5R7ltUL4DTQ
RKdVGLOFIT8Z+pCPrdiuK9M5eqbxWkukrkOCUTXFctJFJyZ52lFgNwHz+Cbrfbuvle8PRvVZzXjR
JT4t5D37onAL8makM6eiQils1s1/JreVXdJd5fe6UP76Rs0sZd9EZDs5FOeEgXszM1SYOhsLdC3U
ihtQmpYPJawU3rZQ0SYLQZR6zG49BiWSWNecD94QHSVyT1f570LuT2hCrYklEC6YLKvar9ZtUWg8
2nhkaAn0YwgV1Tgx0PoEHLsZ62N8pjaUX/njWOEz7/8gXr9hMubopRrKy7KLkcXfUrlP+wdcIfKS
tqfCECh2hIF3r4AM9ycfp//HmrHM1vP9TfVk0hNYmJI5AqUUX2t7sJDjjEVmlLpmYb1LsUNt3Q1l
ZhL2ccFVlVAhhyGV5rKEP4TMWfqckvRIf8rmf4Zr148AHDR3KedgFg1WEugem/PlJgjFkAizDLtm
UCYi23xx9v+J/QylZosScfqW9E31lvS6NKvYfdA87AwnFH+BTYzpXEZYi25RutgVbXSFabuXTOsT
ZAJvCRECopx9VSxurxaQ1XYDqy+61nc0lam8ROIX6sopG8J1QUHrRjeS/LQ68B7vwwhKm+n0HkfN
MoHuT4+4ixGMQic4Cdmobnd/Xf5y29HGlIbgXni6JZJLLK9/qUNL7sMS75jUJThOC509Pz8YQyKl
RLcZJEnde9t7YN5o0J2QI7Dlvtqd9cYSLdKYBOH76IsZZ60mawADVGsoZcBb2GbCUP9SDv1NSJ41
TlRcjWCZjhg+D9I+uAqpBaKriTD+R6ZFWMRTkvuATCPcJ0cDyittckydcUBZbhVZmChUpUhogYz2
zwe5YvYRKhT34X9O+/VV+QfnigCFMLoqGEgSCqEPR4vgn3S2aGVjgI4cuQ+7SOxAt1TX3sINxGmT
HAdfo2hKoJrwTb1eXFuHWI8AEsFC/0c2YGFwpw4OiYGZspuZbhBd5qkz11mCe3ogdI0sh34ywLx+
5fvE5SSfHBkwGB+rTAWssWRRZlIeE1k3AHmRcaXt2bxGwOKkrTMUlHoKNCTgF7Ez/aqIYrRRPKZa
zWRA8L/HEe/hlFLoPg76B81volNoo793qBePE7S0uYJQkEzogUxi3KC+z9jjMbZTdSr3+f+2vZbp
X3TVjjRj8mYyBXARwRPvSWxcl4eCLpvRRkRqQ+sKsV7j92BS5EsM/aKEx/wdMeV6OYvj/vSu3Hly
xqn5B0NuYzSkmdJkWBx8woWW/8IJJ84Nrph4RD1ypg4mIcyle8LM5a1Hul3kbmWJGIJooOyquscC
XeiGnTI/Ai1sYyKzg9XiDfLdv3qBUv4DZNrlcPRNkLvyKSTqQJxBPOycvc5gr8AYwuE2FLu6zW5x
yCIrnYjy+P4W1LbcVqTT2GSRyIjZtUWCqOVGt4M7dbslJwZyn2olSwufZTCoIzGr+NEBS2P7+o/M
0KTejlQnykvk19gungZYjl9WHmUZtDhe6VLXCDrBIFuypWY0ch7FmhJaQPCw6DEJ3EuN/nEyArlh
N+2LycHvJ2X4hB4CyuieziR2qo2rW63ZaT1w27p7LDp6/38+oohOjotO+uq6mbQyEdzhcpO54Eyc
iwr4QSu+B1cuYUFg9xTNqRW+mPtA1yk13Z0KL0qpI+YJFIBFcvGMpn0/Gm585EoAQyeMYgFuuS7I
9jaoY5dE8SK+upfAQ2Mw6DggD0vV4fbIud6Y4G8aDP2gRyIlvjfnwnzNgm9OQbXT9E5kNoaa7kWK
b8T0pK6dgErpJsIoTtnFOcuOCS9LE2pEY6FC1i5XvE/fHdMBXEGkYfQUjChZiBfQi0zRtUWETOnh
pZy4FXIsIgusfuGKApTsqbyU/NBX9CFLgpzCxFuFsNco2sUI4t7RypP098INuCfWn7/HTMtjqtsx
F3MAijHVjWCJ2QfBqGFYEl848dVkTANBMC8r7A2GFgro1skWyaTSVyFI861WPgOwvpJOhSinPHSu
X3dNl2F8yGZom9BulhkjxHpqfuU53RdzpqTSsObfnMaE0AlNKXOzkXLnUaST7sYoBXxt85eIooNe
Dt8iAyErLS9BH8jI/CwUtVTVETAh2lp7MMuJabtXAHbhs8ycx7Hz3yPq03nwCJK2tA6kSoZ58Eux
+qfL/hCuQCWBqYLnLOv/4SR93YZELjRbipRK86dVmKDXMVRV/yfnwBfk5a7PRhK+Og8b54e5CjHq
ZFmatFMlht5Q+f1/FbO49AsXYfc+n6xqm8NfLxyJDiiqN0BVZ4hggw1hEAJEz7k5FpxgHz1Q+9uG
hwgAY5K8JsVLokvLon7h2h2XpL/JBaTLGXRGve2g6Ijfvtwv7npX/XVWH2Zfm/aim2yiuC5tC1rY
qOyO21OoSBJ1iri1IH0eDNFak/AO6xDLw4+Hcv6ZKsenP1dPd9pEpnvC1YwIItO3j9sWOFWlEw1Z
mq+Xwxfyv7aLP7rKRqkEUiPt+UYrskFpcuVEV9RdfgtMvbsn2Q9o+N2g/NZSx2pxiGCAwM4DmHoz
Y6xipRmzcgo30G4ZoPQSG7/GWIejm6FZ3duP8qwZCRVV1DZlXHSE15TofLAs2rTBY2yWRGTvkMF/
JDA4cVLKXEw2e8Ro+eB0PGipC9KnuMrzKF6h2QGXAUkxsWv8tKmqdEWT0b9ixJ+GTVHdd4vK8j3V
oSnLnmpnMkx8a75mF1mU6LaR5PFMdEIfsWpbrnBs+QTtI3+cg52jhmzQCq+3U+DoMxmEyfT9OTiq
T6pl5yPuXdU9wl2rPEKbVxFavT/ULwFJoMaVHHi1tu5Tc5YnHV4y42zRqP55Ith8GDZP+b1p47Z8
NPCjGSpBFV5tOFBOegjwl5bdcdZldfOuQAj6ZqinNBaVjkeECMtulh/ygYUpRiSg9CfEjigeUUWo
UeSC5oFuKjMFKdHDiZap231X3AXzEGw//2OO5+st6m0LLKMmgUWjchoIb/b2pvLcr6S78m0VtdHK
VFaBt5fbh+8CWKneWnoqClW0W0MeOvzhXqP15icKrh3JXNlkK/h8qqjnem41g7GIgb7wac3rhet2
ceaY3DvuxFV1/P54bbCXeJuHReYt2eCHH9k+4PT7VRYt+No3pYmC4XZoe6FxOXk+CxkvNkRXxO9P
+JrTqFr1ZCAAgdCS4CBiljD31fu5/vFfKIdFepeSBYW4DE6y7eMbAauZM//itSqdPDaAXY3cRKyI
LoX7xLK1BmJA/L1rEPTnbTLzdq+ejbV+zEZN6V67IHdLzsLjYI/Fnr2styhKGe3d2RzU2JdDWDwW
yZrDhKsqBHKFYzjeRpIQ9iLxUobfWY5Zjm7Izw8xvsPowTzil+Iasd8WO7ppzdmQp1K22Chw55Yh
2Ev5dV/W8hJ+JQkZRD+fm/JewdzxVmWLmOtM5WSEjj1WpZp3tMCcQTeXM2bccBb28iMM/yeUkdqX
DqRtVU/0vcgHsjBPhCI8+tkenoJFovTiBPTnTQq78CYGEeGuLkp8/mzZ4HZEb+H6WWnZQyLK+sCD
89k9aqHOHtRmdx7c8CPSD+ZBRmskxEKsivDXMionAGWF7OSQkaOuTeMkHZIm7kgvEp6intj91/Pg
kZSY2651/ED+wXBhoX0W8RwkegvPRGR4QsGbY6u4wUDJViJPrmzjcLdAR8AU4II0JmSBTCW93rUC
hvFqtk46+P6b6NRXvBvy+BxgBCQgExrlgpyMQtH4N8xkhUCCq6sTGJgPTQ==
`protect end_protected
